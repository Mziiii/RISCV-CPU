// `include "config.v"

// module alu (
//     input wire clk,
//     input wire rst,
//     input wire rdy,

//     // request(add-inst) from alu_rs
//     input wire alu_en_i,
//     input wire [`OpBus] opcode_i,
//     input wire [`DataBus] rs1_i,
//     input wire [`DataBus] rs2_i,
//     input wire [`] ;


//     input wire [`DataBus] 
// );

// always @(*) begin
    
// end

// always @(posedge clk) begin
    
// end
    
// endmodule