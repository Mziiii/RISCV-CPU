// `include "config.v"

// module alu_rs (
//     input wire clk,
//     input wire rst,
//     input wire rdy,

//     input wire clear,

//     //dispatch 
//     input wire dp_en_i,
//     input wire [`OpBus] op_i,
//     input wire [`ImmBus] imm_i,
//     input wire [`AddrBus] pc_i,
//     input wire [`TagBus] des_i,

//     input wire 
// );
    
// endmodule
